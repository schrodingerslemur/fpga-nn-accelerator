// Common parameters
`ifndef DEFS_SVH
`define DEFS_SVH


`define DATA_WIDTH 16
`define ACC_WIDTH 32


`endif